// wpa2.v

// Generated using ACDS version 15.1 185

`timescale 1 ps / 1 ps
module wpa2 (
		output wire [7:0]  address_export,                  //                  address.export
		input  wire        altpll_areset_conduit_export,    //    altpll_areset_conduit.export
		output wire        altpll_locked_conduit_export,    //    altpll_locked_conduit.export
		output wire        altpll_phasedone_conduit_export, // altpll_phasedone_conduit.export
		input  wire        clk_clk,                         //                      clk.clk
		inout  wire [7:0]  control_export,                  //                  control.export
		output wire [11:0] ram_wire_addr,                   //                 ram_wire.addr
		output wire [1:0]  ram_wire_ba,                     //                         .ba
		output wire        ram_wire_cas_n,                  //                         .cas_n
		output wire        ram_wire_cke,                    //                         .cke
		output wire        ram_wire_cs_n,                   //                         .cs_n
		inout  wire [15:0] ram_wire_dq,                     //                         .dq
		output wire [1:0]  ram_wire_dqm,                    //                         .dqm
		output wire        ram_wire_ras_n,                  //                         .ras_n
		output wire        ram_wire_we_n,                   //                         .we_n
		input  wire [31:0] read_export,                     //                     read.export
		input  wire        reset_reset_n,                   //                    reset.reset_n
		output wire [31:0] write_export                     //                    write.export
	);

	wire         altpll_c0_clk;                                             // altpll:c0 -> [irq_mapper:clk, jtag_uart:clk, mm_interconnect_0:altpll_c0_clk, nios2_e:clk, onchip_memory:clk, pio_address:clk, pio_control:clk, pio_read_data:clk, pio_write_data:clk, rst_controller_001:clk, sdram_controller:clk]
	wire  [31:0] nios2_e_data_master_readdata;                              // mm_interconnect_0:nios2_e_data_master_readdata -> nios2_e:d_readdata
	wire         nios2_e_data_master_waitrequest;                           // mm_interconnect_0:nios2_e_data_master_waitrequest -> nios2_e:d_waitrequest
	wire         nios2_e_data_master_debugaccess;                           // nios2_e:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_e_data_master_debugaccess
	wire  [24:0] nios2_e_data_master_address;                               // nios2_e:d_address -> mm_interconnect_0:nios2_e_data_master_address
	wire   [3:0] nios2_e_data_master_byteenable;                            // nios2_e:d_byteenable -> mm_interconnect_0:nios2_e_data_master_byteenable
	wire         nios2_e_data_master_read;                                  // nios2_e:d_read -> mm_interconnect_0:nios2_e_data_master_read
	wire         nios2_e_data_master_write;                                 // nios2_e:d_write -> mm_interconnect_0:nios2_e_data_master_write
	wire  [31:0] nios2_e_data_master_writedata;                             // nios2_e:d_writedata -> mm_interconnect_0:nios2_e_data_master_writedata
	wire  [31:0] nios2_e_instruction_master_readdata;                       // mm_interconnect_0:nios2_e_instruction_master_readdata -> nios2_e:i_readdata
	wire         nios2_e_instruction_master_waitrequest;                    // mm_interconnect_0:nios2_e_instruction_master_waitrequest -> nios2_e:i_waitrequest
	wire  [24:0] nios2_e_instruction_master_address;                        // nios2_e:i_address -> mm_interconnect_0:nios2_e_instruction_master_address
	wire         nios2_e_instruction_master_read;                           // nios2_e:i_read -> mm_interconnect_0:nios2_e_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_nios2_e_debug_mem_slave_readdata;        // nios2_e:debug_mem_slave_readdata -> mm_interconnect_0:nios2_e_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_e_debug_mem_slave_waitrequest;     // nios2_e:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_e_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_e_debug_mem_slave_debugaccess;     // mm_interconnect_0:nios2_e_debug_mem_slave_debugaccess -> nios2_e:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_e_debug_mem_slave_address;         // mm_interconnect_0:nios2_e_debug_mem_slave_address -> nios2_e:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_e_debug_mem_slave_read;            // mm_interconnect_0:nios2_e_debug_mem_slave_read -> nios2_e:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_e_debug_mem_slave_byteenable;      // mm_interconnect_0:nios2_e_debug_mem_slave_byteenable -> nios2_e:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_e_debug_mem_slave_write;           // mm_interconnect_0:nios2_e_debug_mem_slave_write -> nios2_e:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_e_debug_mem_slave_writedata;       // mm_interconnect_0:nios2_e_debug_mem_slave_writedata -> nios2_e:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_altpll_pll_slave_readdata;               // altpll:readdata -> mm_interconnect_0:altpll_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_altpll_pll_slave_address;                // mm_interconnect_0:altpll_pll_slave_address -> altpll:address
	wire         mm_interconnect_0_altpll_pll_slave_read;                   // mm_interconnect_0:altpll_pll_slave_read -> altpll:read
	wire         mm_interconnect_0_altpll_pll_slave_write;                  // mm_interconnect_0:altpll_pll_slave_write -> altpll:write
	wire  [31:0] mm_interconnect_0_altpll_pll_slave_writedata;              // mm_interconnect_0:altpll_pll_slave_writedata -> altpll:writedata
	wire         mm_interconnect_0_onchip_memory_s1_chipselect;             // mm_interconnect_0:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_readdata;               // onchip_memory:readdata -> mm_interconnect_0:onchip_memory_s1_readdata
	wire  [12:0] mm_interconnect_0_onchip_memory_s1_address;                // mm_interconnect_0:onchip_memory_s1_address -> onchip_memory:address
	wire   [3:0] mm_interconnect_0_onchip_memory_s1_byteenable;             // mm_interconnect_0:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	wire         mm_interconnect_0_onchip_memory_s1_write;                  // mm_interconnect_0:onchip_memory_s1_write -> onchip_memory:write
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_writedata;              // mm_interconnect_0:onchip_memory_s1_writedata -> onchip_memory:writedata
	wire         mm_interconnect_0_onchip_memory_s1_clken;                  // mm_interconnect_0:onchip_memory_s1_clken -> onchip_memory:clken
	wire         mm_interconnect_0_pio_address_s1_chipselect;               // mm_interconnect_0:pio_address_s1_chipselect -> pio_address:chipselect
	wire  [31:0] mm_interconnect_0_pio_address_s1_readdata;                 // pio_address:readdata -> mm_interconnect_0:pio_address_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_address_s1_address;                  // mm_interconnect_0:pio_address_s1_address -> pio_address:address
	wire         mm_interconnect_0_pio_address_s1_write;                    // mm_interconnect_0:pio_address_s1_write -> pio_address:write_n
	wire  [31:0] mm_interconnect_0_pio_address_s1_writedata;                // mm_interconnect_0:pio_address_s1_writedata -> pio_address:writedata
	wire         mm_interconnect_0_pio_write_data_s1_chipselect;            // mm_interconnect_0:pio_write_data_s1_chipselect -> pio_write_data:chipselect
	wire  [31:0] mm_interconnect_0_pio_write_data_s1_readdata;              // pio_write_data:readdata -> mm_interconnect_0:pio_write_data_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_write_data_s1_address;               // mm_interconnect_0:pio_write_data_s1_address -> pio_write_data:address
	wire         mm_interconnect_0_pio_write_data_s1_write;                 // mm_interconnect_0:pio_write_data_s1_write -> pio_write_data:write_n
	wire  [31:0] mm_interconnect_0_pio_write_data_s1_writedata;             // mm_interconnect_0:pio_write_data_s1_writedata -> pio_write_data:writedata
	wire  [31:0] mm_interconnect_0_pio_read_data_s1_readdata;               // pio_read_data:readdata -> mm_interconnect_0:pio_read_data_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_read_data_s1_address;                // mm_interconnect_0:pio_read_data_s1_address -> pio_read_data:address
	wire         mm_interconnect_0_pio_control_s1_chipselect;               // mm_interconnect_0:pio_control_s1_chipselect -> pio_control:chipselect
	wire  [31:0] mm_interconnect_0_pio_control_s1_readdata;                 // pio_control:readdata -> mm_interconnect_0:pio_control_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_control_s1_address;                  // mm_interconnect_0:pio_control_s1_address -> pio_control:address
	wire         mm_interconnect_0_pio_control_s1_write;                    // mm_interconnect_0:pio_control_s1_write -> pio_control:write_n
	wire  [31:0] mm_interconnect_0_pio_control_s1_writedata;                // mm_interconnect_0:pio_control_s1_writedata -> pio_control:writedata
	wire         mm_interconnect_0_sdram_controller_s1_chipselect;          // mm_interconnect_0:sdram_controller_s1_chipselect -> sdram_controller:az_cs
	wire  [15:0] mm_interconnect_0_sdram_controller_s1_readdata;            // sdram_controller:za_data -> mm_interconnect_0:sdram_controller_s1_readdata
	wire         mm_interconnect_0_sdram_controller_s1_waitrequest;         // sdram_controller:za_waitrequest -> mm_interconnect_0:sdram_controller_s1_waitrequest
	wire  [21:0] mm_interconnect_0_sdram_controller_s1_address;             // mm_interconnect_0:sdram_controller_s1_address -> sdram_controller:az_addr
	wire         mm_interconnect_0_sdram_controller_s1_read;                // mm_interconnect_0:sdram_controller_s1_read -> sdram_controller:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_controller_s1_byteenable;          // mm_interconnect_0:sdram_controller_s1_byteenable -> sdram_controller:az_be_n
	wire         mm_interconnect_0_sdram_controller_s1_readdatavalid;       // sdram_controller:za_valid -> mm_interconnect_0:sdram_controller_s1_readdatavalid
	wire         mm_interconnect_0_sdram_controller_s1_write;               // mm_interconnect_0:sdram_controller_s1_write -> sdram_controller:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_controller_s1_writedata;           // mm_interconnect_0:sdram_controller_s1_writedata -> sdram_controller:az_data
	wire         irq_mapper_receiver0_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_e_irq_irq;                                           // irq_mapper:sender_irq -> nios2_e:irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [altpll:reset, mm_interconnect_0:altpll_inclk_interface_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset;                        // rst_controller_001:reset_out -> [irq_mapper:reset, jtag_uart:rst_n, mm_interconnect_0:nios2_e_reset_reset_bridge_in_reset_reset, nios2_e:reset_n, onchip_memory:reset, pio_address:reset_n, pio_control:reset_n, pio_read_data:reset_n, pio_write_data:reset_n, rst_translator:in_reset, sdram_controller:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                    // rst_controller_001:reset_req -> [nios2_e:reset_req, onchip_memory:reset_req, rst_translator:reset_req_in]

	wpa2_altpll altpll (
		.clk       (clk_clk),                                      //       inclk_interface.clk
		.reset     (rst_controller_reset_out_reset),               // inclk_interface_reset.reset
		.read      (mm_interconnect_0_altpll_pll_slave_read),      //             pll_slave.read
		.write     (mm_interconnect_0_altpll_pll_slave_write),     //                      .write
		.address   (mm_interconnect_0_altpll_pll_slave_address),   //                      .address
		.readdata  (mm_interconnect_0_altpll_pll_slave_readdata),  //                      .readdata
		.writedata (mm_interconnect_0_altpll_pll_slave_writedata), //                      .writedata
		.c0        (altpll_c0_clk),                                //                    c0.clk
		.areset    (altpll_areset_conduit_export),                 //        areset_conduit.export
		.locked    (altpll_locked_conduit_export),                 //        locked_conduit.export
		.phasedone (altpll_phasedone_conduit_export)               //     phasedone_conduit.export
	);

	wpa2_jtag_uart jtag_uart (
		.clk            (altpll_c0_clk),                                             //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	wpa2_nios2_e nios2_e (
		.clk                                 (altpll_c0_clk),                                         //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                   //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),                //                          .reset_req
		.d_address                           (nios2_e_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_e_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_e_data_master_read),                              //                          .read
		.d_readdata                          (nios2_e_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_e_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_e_data_master_write),                             //                          .write
		.d_writedata                         (nios2_e_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_e_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_e_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_e_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_e_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_e_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_e_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                      //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_e_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_e_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_e_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_e_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_e_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_e_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_e_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_e_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                       // custom_instruction_master.readra
	);

	wpa2_onchip_memory onchip_memory (
		.clk        (altpll_c0_clk),                                 //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),            // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req)         //       .reset_req
	);

	wpa2_pio_address pio_address (
		.clk        (altpll_c0_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_pio_address_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_address_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_address_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_address_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_address_s1_readdata),   //                    .readdata
		.out_port   (address_export)                               // external_connection.export
	);

	wpa2_pio_control pio_control (
		.clk        (altpll_c0_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_pio_control_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_control_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_control_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_control_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_control_s1_readdata),   //                    .readdata
		.bidir_port (control_export)                               // external_connection.export
	);

	wpa2_pio_read_data pio_read_data (
		.clk      (altpll_c0_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),         //               reset.reset_n
		.address  (mm_interconnect_0_pio_read_data_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_read_data_s1_readdata), //                    .readdata
		.in_port  (read_export)                                  // external_connection.export
	);

	wpa2_pio_write_data pio_write_data (
		.clk        (altpll_c0_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_pio_write_data_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_write_data_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_write_data_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_write_data_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_write_data_s1_readdata),   //                    .readdata
		.out_port   (write_export)                                    // external_connection.export
	);

	wpa2_sdram_controller sdram_controller (
		.clk            (altpll_c0_clk),                                       //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),                 // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_controller_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_controller_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_controller_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_controller_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_controller_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_controller_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_controller_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_controller_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_controller_s1_waitrequest),   //      .waitrequest
		.zs_addr        (ram_wire_addr),                                       //  wire.export
		.zs_ba          (ram_wire_ba),                                         //      .export
		.zs_cas_n       (ram_wire_cas_n),                                      //      .export
		.zs_cke         (ram_wire_cke),                                        //      .export
		.zs_cs_n        (ram_wire_cs_n),                                       //      .export
		.zs_dq          (ram_wire_dq),                                         //      .export
		.zs_dqm         (ram_wire_dqm),                                        //      .export
		.zs_ras_n       (ram_wire_ras_n),                                      //      .export
		.zs_we_n        (ram_wire_we_n)                                        //      .export
	);

	wpa2_mm_interconnect_0 mm_interconnect_0 (
		.altpll_c0_clk                                            (altpll_c0_clk),                                             //                                          altpll_c0.clk
		.clk_48_clk_clk                                           (clk_clk),                                                   //                                         clk_48_clk.clk
		.altpll_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // altpll_inclk_interface_reset_reset_bridge_in_reset.reset
		.nios2_e_reset_reset_bridge_in_reset_reset                (rst_controller_001_reset_out_reset),                        //                nios2_e_reset_reset_bridge_in_reset.reset
		.nios2_e_data_master_address                              (nios2_e_data_master_address),                               //                                nios2_e_data_master.address
		.nios2_e_data_master_waitrequest                          (nios2_e_data_master_waitrequest),                           //                                                   .waitrequest
		.nios2_e_data_master_byteenable                           (nios2_e_data_master_byteenable),                            //                                                   .byteenable
		.nios2_e_data_master_read                                 (nios2_e_data_master_read),                                  //                                                   .read
		.nios2_e_data_master_readdata                             (nios2_e_data_master_readdata),                              //                                                   .readdata
		.nios2_e_data_master_write                                (nios2_e_data_master_write),                                 //                                                   .write
		.nios2_e_data_master_writedata                            (nios2_e_data_master_writedata),                             //                                                   .writedata
		.nios2_e_data_master_debugaccess                          (nios2_e_data_master_debugaccess),                           //                                                   .debugaccess
		.nios2_e_instruction_master_address                       (nios2_e_instruction_master_address),                        //                         nios2_e_instruction_master.address
		.nios2_e_instruction_master_waitrequest                   (nios2_e_instruction_master_waitrequest),                    //                                                   .waitrequest
		.nios2_e_instruction_master_read                          (nios2_e_instruction_master_read),                           //                                                   .read
		.nios2_e_instruction_master_readdata                      (nios2_e_instruction_master_readdata),                       //                                                   .readdata
		.altpll_pll_slave_address                                 (mm_interconnect_0_altpll_pll_slave_address),                //                                   altpll_pll_slave.address
		.altpll_pll_slave_write                                   (mm_interconnect_0_altpll_pll_slave_write),                  //                                                   .write
		.altpll_pll_slave_read                                    (mm_interconnect_0_altpll_pll_slave_read),                   //                                                   .read
		.altpll_pll_slave_readdata                                (mm_interconnect_0_altpll_pll_slave_readdata),               //                                                   .readdata
		.altpll_pll_slave_writedata                               (mm_interconnect_0_altpll_pll_slave_writedata),              //                                                   .writedata
		.jtag_uart_avalon_jtag_slave_address                      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                        jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                                   .write
		.jtag_uart_avalon_jtag_slave_read                         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                                   .read
		.jtag_uart_avalon_jtag_slave_readdata                     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                                   .readdata
		.jtag_uart_avalon_jtag_slave_writedata                    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                                   .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                                   .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                                   .chipselect
		.nios2_e_debug_mem_slave_address                          (mm_interconnect_0_nios2_e_debug_mem_slave_address),         //                            nios2_e_debug_mem_slave.address
		.nios2_e_debug_mem_slave_write                            (mm_interconnect_0_nios2_e_debug_mem_slave_write),           //                                                   .write
		.nios2_e_debug_mem_slave_read                             (mm_interconnect_0_nios2_e_debug_mem_slave_read),            //                                                   .read
		.nios2_e_debug_mem_slave_readdata                         (mm_interconnect_0_nios2_e_debug_mem_slave_readdata),        //                                                   .readdata
		.nios2_e_debug_mem_slave_writedata                        (mm_interconnect_0_nios2_e_debug_mem_slave_writedata),       //                                                   .writedata
		.nios2_e_debug_mem_slave_byteenable                       (mm_interconnect_0_nios2_e_debug_mem_slave_byteenable),      //                                                   .byteenable
		.nios2_e_debug_mem_slave_waitrequest                      (mm_interconnect_0_nios2_e_debug_mem_slave_waitrequest),     //                                                   .waitrequest
		.nios2_e_debug_mem_slave_debugaccess                      (mm_interconnect_0_nios2_e_debug_mem_slave_debugaccess),     //                                                   .debugaccess
		.onchip_memory_s1_address                                 (mm_interconnect_0_onchip_memory_s1_address),                //                                   onchip_memory_s1.address
		.onchip_memory_s1_write                                   (mm_interconnect_0_onchip_memory_s1_write),                  //                                                   .write
		.onchip_memory_s1_readdata                                (mm_interconnect_0_onchip_memory_s1_readdata),               //                                                   .readdata
		.onchip_memory_s1_writedata                               (mm_interconnect_0_onchip_memory_s1_writedata),              //                                                   .writedata
		.onchip_memory_s1_byteenable                              (mm_interconnect_0_onchip_memory_s1_byteenable),             //                                                   .byteenable
		.onchip_memory_s1_chipselect                              (mm_interconnect_0_onchip_memory_s1_chipselect),             //                                                   .chipselect
		.onchip_memory_s1_clken                                   (mm_interconnect_0_onchip_memory_s1_clken),                  //                                                   .clken
		.pio_address_s1_address                                   (mm_interconnect_0_pio_address_s1_address),                  //                                     pio_address_s1.address
		.pio_address_s1_write                                     (mm_interconnect_0_pio_address_s1_write),                    //                                                   .write
		.pio_address_s1_readdata                                  (mm_interconnect_0_pio_address_s1_readdata),                 //                                                   .readdata
		.pio_address_s1_writedata                                 (mm_interconnect_0_pio_address_s1_writedata),                //                                                   .writedata
		.pio_address_s1_chipselect                                (mm_interconnect_0_pio_address_s1_chipselect),               //                                                   .chipselect
		.pio_control_s1_address                                   (mm_interconnect_0_pio_control_s1_address),                  //                                     pio_control_s1.address
		.pio_control_s1_write                                     (mm_interconnect_0_pio_control_s1_write),                    //                                                   .write
		.pio_control_s1_readdata                                  (mm_interconnect_0_pio_control_s1_readdata),                 //                                                   .readdata
		.pio_control_s1_writedata                                 (mm_interconnect_0_pio_control_s1_writedata),                //                                                   .writedata
		.pio_control_s1_chipselect                                (mm_interconnect_0_pio_control_s1_chipselect),               //                                                   .chipselect
		.pio_read_data_s1_address                                 (mm_interconnect_0_pio_read_data_s1_address),                //                                   pio_read_data_s1.address
		.pio_read_data_s1_readdata                                (mm_interconnect_0_pio_read_data_s1_readdata),               //                                                   .readdata
		.pio_write_data_s1_address                                (mm_interconnect_0_pio_write_data_s1_address),               //                                  pio_write_data_s1.address
		.pio_write_data_s1_write                                  (mm_interconnect_0_pio_write_data_s1_write),                 //                                                   .write
		.pio_write_data_s1_readdata                               (mm_interconnect_0_pio_write_data_s1_readdata),              //                                                   .readdata
		.pio_write_data_s1_writedata                              (mm_interconnect_0_pio_write_data_s1_writedata),             //                                                   .writedata
		.pio_write_data_s1_chipselect                             (mm_interconnect_0_pio_write_data_s1_chipselect),            //                                                   .chipselect
		.sdram_controller_s1_address                              (mm_interconnect_0_sdram_controller_s1_address),             //                                sdram_controller_s1.address
		.sdram_controller_s1_write                                (mm_interconnect_0_sdram_controller_s1_write),               //                                                   .write
		.sdram_controller_s1_read                                 (mm_interconnect_0_sdram_controller_s1_read),                //                                                   .read
		.sdram_controller_s1_readdata                             (mm_interconnect_0_sdram_controller_s1_readdata),            //                                                   .readdata
		.sdram_controller_s1_writedata                            (mm_interconnect_0_sdram_controller_s1_writedata),           //                                                   .writedata
		.sdram_controller_s1_byteenable                           (mm_interconnect_0_sdram_controller_s1_byteenable),          //                                                   .byteenable
		.sdram_controller_s1_readdatavalid                        (mm_interconnect_0_sdram_controller_s1_readdatavalid),       //                                                   .readdatavalid
		.sdram_controller_s1_waitrequest                          (mm_interconnect_0_sdram_controller_s1_waitrequest),         //                                                   .waitrequest
		.sdram_controller_s1_chipselect                           (mm_interconnect_0_sdram_controller_s1_chipselect)           //                                                   .chipselect
	);

	wpa2_irq_mapper irq_mapper (
		.clk           (altpll_c0_clk),                      //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.sender_irq    (nios2_e_irq_irq)                     //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.clk            (altpll_c0_clk),                          //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
